// Implementation of HDMI Spec v1.4a
// By Sameer Puri https://github.com/sameer

module hdmi 
#(
    // Defaults to 640x480 which should be supported by almost if not all HDMI sinks.
    // See README.md or CEA-861-D for enumeration of video id codes.
    // Pixel repetition, interlaced scans and other special output modes are not implemented (yet).
    parameter int VIDEO_ID_CODE = 1
)
(
    input logic clk_pixel_x5,
    input logic clk_pixel,
    input logic clk_audio,
    // synchronous reset back to 0,0
    input logic reset,
    input logic [23:0] rgb,
	 
	 input logic hs_ext,
	 input logic vs_ext,
	 input logic [1:0] mode_ext,

    // These outputs go to your HDMI port
    output logic [2:0] tmds,
    output logic tmds_clock,
	 
	 // These outputs go to your HDMI port, addition
    output logic [2:0] tmds1,
    output logic tmds1_clock,
	 
    
    // All outputs below this line stay inside the FPGA
    // They are used (by you) to pick the color each pixel should have
    // i.e. always_ff @(posedge pixel_clk) rgb <= {8'd0, 8'(cx), 8'(cy)};
    output logic [11:0] cx,
    output logic [10:0] cy,

    // The screen is at the upper left corner of the frame.
    // 0,0 = 0,0 in video
    // the frame includes extra space for sending auxiliary data
    output logic [11:0] frame_width,
    output logic [10:0] frame_height,
    output logic [11:0] screen_width,
    output logic [10:0] screen_height
);

localparam int NUM_CHANNELS = 3;
logic hsync;
logic vsync;

logic [11:0] hsync_porch_start, hsync_porch_size;
logic [10:0] vsync_porch_start, vsync_porch_size;
logic invert;

logic [1:0]  edge_hs, edge_vs;

// See CEA-861-D for more specifics formats described below.
always @ (posedge clk_pixel)
begin
	edge_hs = {edge_hs[0], hs_ext};
	edge_vs = {edge_vs[0], vs_ext};

	case (mode_ext)
	0, 1, 2:
	begin
		frame_width = 896;
		frame_height = 640;
		screen_width = 720;
		screen_height = 576;
		hsync_porch_start = 24;
		hsync_porch_size = 80;
		vsync_porch_start = 7;
		vsync_porch_size = 6;
		invert = 1;
	end
	2:
	begin
		frame_width = 896;
		frame_height = 624;
		screen_width = 720;
		screen_height = 576;
		hsync_porch_start = 24;
		hsync_porch_size = 80;
		vsync_porch_start = 7;
		vsync_porch_size = 6;
		invert = 1;
	end
	3:
	begin
		frame_width = 912;
		frame_height = 622;
		screen_width = 720;
		screen_height = 576;
		hsync_porch_start = 24;
		hsync_porch_size = 80;
		vsync_porch_start = 7;
		vsync_porch_size = 6;
		invert = 1;
	end
	endcase
end

assign hsync = invert ^ (cx >= screen_width + hsync_porch_start && cx < screen_width + hsync_porch_start + hsync_porch_size);
assign vsync = invert ^ (cy >= screen_height + vsync_porch_start && cy < screen_height + vsync_porch_start + vsync_porch_size);



// Wrap-around pixel position counters indicating the pixel to be generated by the user in THIS clock and sent out in the NEXT clock.

logic video_data_period = 0;

logic [2:0] mode = 3'd1;
logic [23:0] video_data = 24'd0;
logic [5:0] control_data = 6'd0;
logic [11:0] data_island_data = 12'd0;

always_ff @(posedge clk_pixel)
begin
	if (reset)
	begin
		cx <= 12'(0);
		cy <= 11'(0);
		  
		video_data_period <= 0;
		  
		mode <= 3'd0;
		video_data <= 24'd0;
		control_data <= 6'd0;
	end
	else
	begin
		if (edge_hs == 2'b01)
			cx <= screen_width + hsync_porch_start;
		else
			cx <= cx == frame_width-1'b1 ? 12'(0) : cx + 1'b1;
			
		if (edge_vs == 2'b01)
			cy <= screen_height + vsync_porch_start;
		else
			cy <= cx == frame_width-1'b1 ? cy == frame_height-1'b1 ? 11'(0) : cy + 1'b1 : cy;
		  
		video_data_period <= cx < screen_width && cy < screen_height;
		
		mode <= video_data_period ? 3'd1 : 3'd0;
		video_data <= rgb;
		control_data <= {4'b0000, {vsync, hsync}}; // ctrl3, ctrl2, ctrl1, ctrl0, vsync, hsync
	end
end



// All logic below relates to the production and output of the 10-bit TMDS code.
logic [9:0] tmds_internal [NUM_CHANNELS-1:0];
genvar i;
generate
    // TMDS code production.
	for (i = 0; i < NUM_CHANNELS; i++)
	begin: tmds_gen
		tmds_channel #(.CN(i)) tmds_channel
		(
			.clk_pixel(clk_pixel),
			.video_data(video_data[i*8+7:i*8]),
			.data_island_data(data_island_data[i*4+3:i*4]),
			.control_data(control_data[i*2+1:i*2]),
			.mode(mode),
			.tmds(tmds_internal[i])
		);
	end
endgenerate



serializer #(.NUM_CHANNELS(NUM_CHANNELS)) 
serializer(
	.clk_pixel(clk_pixel),
	.clk_pixel_x5(clk_pixel_x5),
	.reset(reset),
	.tmds_internal(tmds_internal),
	.tmds(tmds),
	.tmds_clock(tmds_clock)
);

serializer #(.NUM_CHANNELS(NUM_CHANNELS)) 
serializer_1(
	.clk_pixel(clk_pixel),
	.clk_pixel_x5(clk_pixel_x5),
	.reset(reset),
	.tmds_internal(tmds_internal),
	.tmds(tmds1),
	.tmds_clock(tmds1_clock)
);

endmodule
